module test;
   reg cl = 0;
   wire [7:0] alu_out_bus;

   computer Comp(.clk(cl), .alu_out_bus(alu_out_bus));

   initial begin
     $dumpfile("out/dump.vcd");
     $dumpvars(0, test);

     // CAMBIO (a lo huaso): sacamos esta carga manual.
     // Antes: $readmemb("im.dat", Comp.IM.mem);
     // Ahora la 'instruction_memory' se carga solita por dentro, bien arriada.

     // Igual mostramos lo que hay en memoria, pa' que el capataz quede conforme.
     $display("mem[0] = %h", Comp.IM.mem[0]);
     $display("mem[1] = %h", Comp.IM.mem[1]);
     $display("mem[2] = %h", Comp.IM.mem[2]);
     $display("mem[3] = %h", Comp.IM.mem[3]);

     $monitor("At time %t, pc = 0x%h, im = b%b, regA = 0x%h, regB = 0x%h, alu=0x%h (b=0x%h)",
              $time, Comp.pc_out_bus, Comp.im_out_bus, Comp.regA_out_bus, Comp.regB_out_bus, alu_out_bus,
              Comp.im_out_bus[7:0]);

     // Esperamos a que el potro PC llegue a 3 y cerramos la trilla.
     wait (Comp.PC.pc == 3);
     #2;
     $finish;
   end

   // Reloj firme, cada #1 pega un latigazo pa’ avanzar.
   always #1 cl = ~cl;
endmodule
